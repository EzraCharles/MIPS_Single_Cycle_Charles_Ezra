module CP // Priority Encoder (Codificador de prioridad)
#(
	parameter WIDTH = 32,
	parameter SELECTOR = 5
)
(
	input logic 	[SELECTOR-1:0] in,
	output logic 	[WIDTH-1:0] 	out
);

// TODO: how to make this process autonomous?
always_comb
	priority case(in)
		5'b00000	:	out = 32'b00000000_00000000_00000000_00000000;
		5'b00001	:	out = 32'b00000000_00000000_00000000_00000010;
		5'b00010	:	out = 32'b00000000_00000000_00000000_00000100;
		5'b00011	:	out = 32'b00000000_00000000_00000000_00001000;
		5'b00100	:	out = 32'b00000000_00000000_00000000_00010000;
		5'b00101	:	out = 32'b00000000_00000000_00000000_00100000;
		5'b00110	:	out = 32'b00000000_00000000_00000000_01000000;
		5'b00111	:	out = 32'b00000000_00000000_00000000_10000000;
		5'b01000	:	out = 32'b00000000_00000000_00000001_00000000;
		5'b01001	:	out = 32'b00000000_00000000_00000010_00000000;
		5'b01010	:	out = 32'b00000000_00000000_00000100_00000000;
		5'b01011	:	out = 32'b00000000_00000000_00001000_00000000;
		5'b01100	:	out = 32'b00000000_00000000_00010000_00000000;
		5'b01101	:	out = 32'b00000000_00000000_00100000_00000000;
		5'b01110	:	out = 32'b00000000_00000000_01000000_00000000;
		5'b01111	:	out = 32'b00000000_00000000_10000000_00000000;
		5'b10000	:	out = 32'b00000000_00000001_00000000_00000000;
		5'b10001	:	out = 32'b00000000_00000010_00000000_00000000;
		5'b10010	:	out = 32'b00000000_00000100_00000000_00000000;
		5'b10011	:	out = 32'b00000000_00001000_00000000_00000000;
		5'b10100	:	out = 32'b00000000_00010000_00000000_00000000;
		5'b10101	:	out = 32'b00000000_00100000_00000000_00000000;
		5'b10110	:	out = 32'b00000000_01000000_00000000_00000000;
		5'b10111	:	out = 32'b00000000_10000000_00000000_00000000;
		5'b11000	:	out = 32'b00000001_00000000_00000000_00000000;
		5'b11001	:	out = 32'b00000010_00000000_00000000_00000000;
		5'b11010	:	out = 32'b00000100_00000000_00000000_00000000;
		5'b11011	:	out = 32'b00001000_00000000_00000000_00000000;
		5'b11100	:	out = 32'b00010000_00000000_00000000_00000000;
		5'b11101	:	out = 32'b00100000_00000000_00000000_00000000;
		5'b11110	:	out = 32'b01000000_00000000_00000000_00000000;
		5'b11111	:	out = 32'b10000000_00000000_00000000_00000000;
	endcase
	
endmodule
